.global VDD VSS

.subckt TOP A C D
X0 A C B E DINV
X1 E D INVX1
.ends 

.subckt DINV A<1> A<2> B<1> B<2>
XA A<1> B<1> INVX1
XB A<2> B<2> INVX1
.ends

.subckt INVX1 A Z
M0 Z A VSS VSS NMOS W=0.95U L=0.25U
M1 Z A VDD VDD PMOS W=1.5U L=0.25U
.ends 
